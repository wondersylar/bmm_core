  );

  const logic [0:1023] [31:0] mem = {
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h0100006F,
    32'h0100006F,
    32'h0080006F,
    32'h0040006F,
    32'h0000006F,
    32'h30047073,
    32'h00000093,
    32'h00008113,
    32'h00008193,
    32'h00008213,
    32'h00008293,
    32'h00008313,
    32'h00008393,
    32'h00008413,
    32'h00008493,
    32'h00008513,
    32'h00008593,
    32'h00008613,
    32'h00008693,
    32'h00008713,
    32'h00008793,
    32'h00008813,
    32'h00008893,
    32'h00008913,
    32'h00008993,
    32'h00008A13,
    32'h00008A93,
    32'h00008B13,
    32'h00008B93,
    32'h00008C13,
    32'h00008C93,
    32'h00008D13,
    32'h00008D93,
    32'h00008E13,
    32'h00008E93,
    32'h00008F13,
    32'h00008F93,
    32'h00100117,
    32'hCF010113,
    32'h000F8D17,
    32'hEE8D0D13,
    32'h000F8D97,
    32'hEE0D8D93,
    32'h01BD5863,
    32'h000D2023,
    32'h004D0D13,
    32'hFFADDCE3,
    32'h000F8D17,
    32'hEC8D0D13,
    32'h000F8D97,
    32'hEC0D8D93,
    32'h00001C97,
    32'hC28C8C93,
    32'h01BD5C63,
    32'h000CAC03,
    32'h018D2023,
    32'h004D0D13,
    32'h004C8C93,
    32'hFFBD48E3,
    32'h00000513,
    32'h00000593,
    32'h004000EF,
    32'h45957131,
    32'hDF064501,
    32'hDB26DD22,
    32'hD74ED94A,
    32'hD356D552,
    32'hCF5ED15A,
    32'hCB66CD62,
    32'hC76EC96A,
    32'h714000EF,
    32'h05136525,
    32'h00EFC6E5,
    32'h05137660,
    32'h00EF0200,
    32'h05137AE0,
    32'h00EF0200,
    32'h440D7A60,
    32'h05134485,
    32'h00EF0300,
    32'h151379A0,
    32'hD5330034,
    32'h051300A4,
    32'h75130305,
    32'h147D0FF5,
    32'h784000EF,
    32'hFFF431E3,
    32'h00EF4529,
    32'h00EF77A0,
    32'h45817960,
    32'h263D4501,
    32'h45014581,
    32'h45012E71,
    32'h842A26B5,
    32'h00108537,
    32'hE0050513,
    32'h22B000EF,
    32'h28040F63,
    32'h05136509,
    32'h25593285,
    32'h27B74711,
    32'hC3D81A10,
    32'h06400513,
    32'h46812DA5,
    32'h45A14601,
    32'h09F00513,
    32'h2E49C002,
    32'h26ED4561,
    32'h45014581,
    32'h458126F1,
    32'h29194501,
    32'h850A45E1,
    32'h842A29B1,
    32'h9537C511,
    32'h05130000,
    32'hA801C945,
    32'h842A2BE1,
    32'h9537C909,
    32'h05130000,
    32'h00EFC9C5,
    32'hC8416AA0,
    32'h9537A051,
    32'h05130000,
    32'h00EFCA45,
    32'h478369A0,
    32'h49030001,
    32'h97130021,
    32'h47830107,
    32'h05130011,
    32'h07A20200,
    32'hE9338FD9,
    32'h00EF0127,
    32'h05136CA0,
    32'h00EF0200,
    32'h448D6C20,
    32'h97934A25,
    32'h57B30034,
    32'hF41300F9,
    32'h57930FF7,
    32'h85130044,
    32'h74630307,
    32'h851300FA,
    32'h00EF0377,
    32'h37B369E0,
    32'h8513F644,
    32'h74630307,
    32'h851300FA,
    32'h14FD0377,
    32'hB6E32561,
    32'h4529FDF4,
    32'h47022541,
    32'h07B7C711,
    32'h17FD0100,
    32'h00F71763,
    32'h00009537,
    32'hCB050513,
    32'h9537AA45,
    32'h05130000,
    32'h2539CB85,
    32'h460146E1,
    32'h450D45A1,
    32'h05132C65,
    32'h26394000,
    32'h45014581,
    32'h45812CC5,
    32'h2E2D4501,
    32'h40000593,
    32'h2EBD850A,
    32'h16051563,
    32'h12632311,
    32'h89371605,
    32'h09130010,
    32'h0A13E009,
    32'h86CA0021,
    32'h07A00613,
    32'h00EF85D2,
    32'h57830C30,
    32'h876307C1,
    32'h953700A7,
    32'h05130000,
    32'hA8F9CC05,
    32'h00009537,
    32'h0513002C,
    32'h2589CC85,
    32'h9537C511,
    32'h05130000,
    32'hA0D9CD85,
    32'h5B0367A5,
    32'h87930181,
    32'hE963D807,
    32'h44810167,
    32'h0C934A81,
    32'h9D370800,
    32'hA8A50000,
    32'h00009537,
    32'hCE050513,
    32'h5703A045,
    32'h00300041,
    32'h00370793,
    32'h86D68389,
    32'h17FD0785,
    32'h0C079763,
    32'hCF8D0513,
    32'h2BA99ABA,
    32'h235D4525,
    32'h0513809D,
    32'h04850200,
    32'h4D8D2B71,
    32'h97934C25,
    32'hD7B3003D,
    32'hF41300F4,
    32'h57930FF7,
    32'h85130044,
    32'h74630307,
    32'h851300FC,
    32'h2BAD0377,
    32'hF64437B3,
    32'h03078513,
    32'h00FC7463,
    32'h03778513,
    32'h239D1DFD,
    32'hFDFDB7E3,
    32'h2BB94529,
    32'h8B9384DE,
    32'hFD630804,
    32'h46E10764,
    32'h008B9613,
    32'h450D45A1,
    32'h05132275,
    32'h24094000,
    32'h45014581,
    32'h05932C15,
    32'h850A4000,
    32'hC5192CA5,
    32'h00009537,
    32'hC9450513,
    32'hA8A129E1,
    32'hC5112ED5,
    32'h00009537,
    32'hC9C50513,
    32'h5783BFC5,
    32'hD7630041,
    32'h953700FC,
    32'h05130000,
    32'hBFF9CE85,
    32'h061386CA,
    32'h85D207A0,
    32'h7A4000EF,
    32'h07C15783,
    32'hF2A787E3,
    32'h00009537,
    32'hCF050513,
    32'h258BB7C1,
    32'hA22B0046,
    32'hB72500B6,
    32'hFD4D2675,
    32'h00009537,
    32'hD2050513,
    32'h2E79A89D,
    32'h9537C511,
    32'h05130000,
    32'h298DC9C5,
    32'h00009537,
    32'hD2850513,
    32'h29D921A5,
    32'h00009537,
    32'hD0850513,
    32'h21E929B1,
    32'h23D14501,
    32'h07B7C91D,
    32'hC7938000,
    32'h953EFEF7,
    32'hE963478D,
    32'h67A500A7,
    32'h8793050A,
    32'hF503D507,
    32'hA02920A7,
    32'h00009537,
    32'hC9050513,
    32'h95372135,
    32'h05130000,
    32'h210DD105,
    32'h2179A001,
    32'h000F4537,
    32'h24050513,
    32'h95372645,
    32'h05130000,
    32'h2129D185,
    32'h77B729A5,
    32'hA4231A10,
    32'h07930007,
    32'h87820800,
    32'h00010001,
    32'hA0010001,
    32'h1A1017B7,
    32'h0007A783,
    32'hFF010113,
    32'h00F12623,
    32'h00100793,
    32'h00C12703,
    32'h00A797B3,
    32'h00059863,
    32'hFFF7C793,
    32'h00E7F7B3,
    32'h0080006F,
    32'h00E7E7B3,
    32'h00F12623,
    32'h00C12703,
    32'h1A1017B7,
    32'h00E7A023,
    32'h01010113,
    32'h00008067,
    32'h1A1017B7,
    32'hFF010113,
    32'h0047A783,
    32'h00F12623,
    32'h00C12783,
    32'h40A7D533,
    32'hFC153533,
    32'h00A12623,
    32'h00C12503,
    32'h01010113,
    32'h00008067,
    32'h1A101737,
    32'h00C70713,
    32'h00100793,
    32'h00072683,
    32'h00A797B3,
    32'h00059863,
    32'hFFF7C513,
    32'h00D577B3,
    32'h0080006F,
    32'h00D7E7B3,
    32'h00F72023,
    32'h00008067,
    32'h02000793,
    32'h40B787B3,
    32'h00F51533,
    32'h1A1027B7,
    32'h00878713,
    32'h00A72023,
    32'h00C78713,
    32'h00C72023,
    32'h00004737,
    32'h00869693,
    32'hF0070713,
    32'h00E6F6B3,
    32'hF265B5B3,
    32'h00B6E5B3,
    32'h01078793,
    32'h00B7A023,
    32'h00008067,
    32'h01059593,
    32'h10055533,
    32'h00A5E5B3,
    32'h1A1027B7,
    32'h00B7AA23,
    32'h00008067,
    32'h1A102737,
    32'h01070713,
    32'h00072783,
    32'hFF010113,
    32'h00F12623,
    32'h00C12783,
    32'h1007D7B3,
    32'h01051513,
    32'h00F56533,
    32'h00A12623,
    32'h00C12783,
    32'h00F72023,
    32'h01010113,
    32'h00008067,
    32'h00100793,
    32'h00858593,
    32'h00001737,
    32'h00B795B3,
    32'h00A79533,
    32'hF0070713,
    32'h00E5F5B3,
    32'hEE853533,
    32'h00A5E533,
    32'h1A1027B7,
    32'h00A7A023,
    32'h00008067,
    32'h1A1027B7,
    32'h0007A783,
    32'hFF010113,
    32'h00F12623,
    32'h00C12503,
    32'h01010113,
    32'h00008067,
    32'h4055D793,
    32'hFC010113,
    32'hE8B7B7B3,
    32'h00F12423,
    32'hF455B7B3,
    32'h03412423,
    32'h02112E23,
    32'h02812C23,
    32'h02912A23,
    32'h03212823,
    32'h03312623,
    32'h03512223,
    32'h03612023,
    32'h01712E23,
    32'h00050A13,
    32'h00078863,
    32'h00812783,
    32'h00178793,
    32'h00F12423,
    32'h4035D593,
    32'h05F5E4B7,
    32'h1A102AB7,
    32'h00010937,
    32'hFA25B433,
    32'h00012623,
    32'h10048493,
    32'h01000B13,
    32'h020A8B93,
    32'hF0090913,
    32'h00FF09B7,
    32'h01010793,
    32'h00C12703,
    32'hFF87A783,
    32'h04F75063,
    32'h000AA783,
    32'h4107D793,
    32'hEE87B7B3,
    32'h02079C63,
    32'h02048063,
    32'h01000513,
    32'h158000EF,
    32'h009B7663,
    32'hFF048493,
    32'hFDDFF06F,
    32'h00000493,
    32'hFD5FF06F,
    32'h80000537,
    32'h00450513,
    32'h0A00006F,
    32'h00000513,
    32'h0980006F,
    32'h000BA783,
    32'h00812703,
    32'hFFF70713,
    32'h00C12683,
    32'h00E6C463,
    32'h02041463,
    32'h0137F733,
    32'h01879613,
    32'h0187D693,
    32'h0127F7B3,
    32'h00D666B3,
    32'h00879793,
    32'h00875713,
    32'h00F6E7B3,
    32'h0180006F,
    32'h00243E63,
    32'h00879713,
    32'h0127F7B3,
    32'hDF073733,
    32'h0087D793,
    32'h00F767B3,
    32'h0240006F,
    32'h02343063,
    32'h0127F6B3,
    32'hEE87B733,
    32'h0137F7B3,
    32'h01071713,
    32'h0107D793,
    32'h00F767B3,
    32'h00F6E7B3,
    32'h00C12703,
    32'h00271713,
    32'h00FA6723,
    32'h00C12783,
    32'h00178793,
    32'h00F12623,
    32'hF1DFF06F,
    32'h03C12083,
    32'h03812403,
    32'h03412483,
    32'h03012903,
    32'h02C12983,
    32'h02812A03,
    32'h02412A83,
    32'h02012B03,
    32'h01C12B83,
    32'h04010113,
    32'h00008067,
    32'hFF010113,
    32'h00812423,
    32'h05F5E437,
    32'h00912223,
    32'h00112623,
    32'h10040413,
    32'h01000493,
    32'hE3DFF0EF,
    32'h10055533,
    32'h02152863,
    32'h02040063,
    32'h01000513,
    32'h03C000EF,
    32'h0084F663,
    32'hFF040413,
    32'hFE1FF06F,
    32'h00000413,
    32'hFD9FF06F,
    32'h80000537,
    32'h00350513,
    32'h0080006F,
    32'h00000513,
    32'h00C12083,
    32'h00812403,
    32'h00412483,
    32'h01010113,
    32'h00008067,
    32'h00150513,
    32'hFFF50513,
    32'h00051463,
    32'h00008067,
    32'h00000013,
    32'hFF1FF06F,
    32'h1A1077B7,
    32'h00478793,
    32'h0007A703,
    32'h0085D613,
    32'hC0174733,
    32'h00E7A023,
    32'h1A1007B7,
    32'h00C78693,
    32'h08300713,
    32'h00E6A023,
    32'h0FF5F593,
    32'h00478713,
    32'h00C72023,
    32'h00B7A42B,
    32'h0A700613,
    32'h00C7A023,
    32'h00300793,
    32'h00F6A023,
    32'h00072783,
    32'h0F07F793,
    32'hC017C7B3,
    32'h00F72023,
    32'h00008067,
    32'h1A1007B7,
    32'h01478793,
    32'h0015468B,
    32'h00068E63,
    32'h0007A703,
    32'h02077713,
    32'hFE070CE3,
    32'h1A100737,
    32'h00D72023,
    32'hFE5FF06F,
    32'h00008067,
    32'h1A100737,
    32'h01470713,
    32'h00072783,
    32'hFC17B7B3,
    32'hFE078CE3,
    32'h1A1007B7,
    32'h0007A503,
    32'h0FF57513,
    32'h00008067,
    32'h1A100737,
    32'h01470713,
    32'h00072783,
    32'h0207F793,
    32'hFE078CE3,
    32'h1A1007B7,
    32'h00A7A023,
    32'h00008067,
    32'h1A100737,
    32'h01470713,
    32'h00072783,
    32'h0407F793,
    32'hFE078CE3,
    32'h00008067,
    32'h1A100537,
    32'h01452503,
    32'hFC153533,
    32'h00008067,
    32'h00B567B3,
    32'hFA27B7B3,
    32'h04079E63,
    32'hFEFF0637,
    32'h80808837,
    32'h00058713,
    32'h00050693,
    32'hEFF60613,
    32'h08080813,
    32'h00070593,
    32'h00068513,
    32'h0005A883,
    32'h0046A78B,
    32'h00470713,
    32'h03179663,
    32'h00C785B3,
    32'hFFF7C793,
    32'h00F5F7B3,
    32'h0107F7B3,
    32'hFC078CE3,
    32'h00000513,
    32'h00008067,
    32'h00074683,
    32'h00158593,
    32'h00F69863,
    32'h0015478B,
    32'h00058713,
    32'hFE0796E3,
    32'h00074503,
    32'h40A78533,
    32'h00008067,
    32'hC4221141,
    32'hC606C226,
    32'h0493842A,
    32'hCC197D00,
    32'hC5093795,
    32'h45333711,
    32'hA8111005,
    32'h7D000513,
    32'hF5633DA1,
    32'h04130084,
    32'hB7D58304,
    32'h2083557D,
    32'h240300C1,
    32'h24830081,
    32'h01410041,
    32'h67A18082,
    32'h060517FD,
    32'h00A7EA63,
    32'hE211167D,
    32'hC78BA031,
    32'h00AB0015,
    32'hBFCD00F5,
    32'h71318082,
    32'hDB26DD22,
    32'h01000437,
    32'h001E84B7,
    32'hD74ED94A,
    32'hDF06D552,
    32'hD15AD356,
    32'hCD62CF5E,
    32'h8A2ACB66,
    32'h48048493,
    32'h09934961,
    32'h04490420,
    32'h3F9D8526,
    32'h04054063,
    32'h0FF57793,
    32'h02F96463,
    32'h00F45733,
    32'hFC173733,
    32'h4985CF11,
    32'h00108AB7,
    32'h4401894E,
    32'h0B134BE1,
    32'h0C130640,
    32'h8A930850,
    32'hA8B1E00A,
    32'h0DF7F793,
    32'hFD3794E3,
    32'h80000537,
    32'hA0ED054D,
    32'h04300513,
    32'hBF5D35B5,
    32'h80AB0405,
    32'h066300AC,
    32'h85260184,
    32'h59E33705,
    32'h4783FE05,
    32'h470300A1,
    32'hC7930091,
    32'hF793FFF7,
    32'h08630FF7,
    32'h455502F7,
    32'h44013581,
    32'h3DFD8526,
    32'h4E630405,
    32'h07130805,
    32'h77930640,
    32'h0A630FF5,
    32'hB96308E4,
    32'h04230417,
    32'h0C9300F1,
    32'h843E0091,
    32'h1AE3BF6D,
    32'h86D6FCE9,
    32'h08000613,
    32'h00B10593,
    32'h207D4501,
    32'h08B14783,
    32'h08C14703,
    32'h97BA07A2,
    32'h1007D7B3,
    32'hFAF519E3,
    32'h09058552,
    32'h08000613,
    32'h00B10593,
    32'h791335DD,
    32'h09850FF9,
    32'h080A0A13,
    32'hBF594519,
    32'h0047BD63,
    32'h33F94519,
    32'h10000793,
    32'hFF634501,
    32'h05370337,
    32'h05458000,
    32'h9B63A815,
    32'h45110177,
    32'h05373B55,
    32'h05498000,
    32'h0405A015,
    32'h01640963,
    32'h359D8526,
    32'hFE054BE3,
    32'h1FE3A039,
    32'h0537F564,
    32'h05518000,
    32'h7793A021,
    32'hB7950FF5,
    32'h0BC12083,
    32'h0B812403,
    32'h0B412483,
    32'h0B012903,
    32'h0AC12983,
    32'h0A812A03,
    32'h0A412A83,
    32'h0A012B03,
    32'h09C12B83,
    32'h09812C03,
    32'h09412C83,
    32'h80826129,
    32'h00160713,
    32'h02065063,
    32'hA8294705,
    32'h0015C78B,
    32'h00855613,
    32'h07868FB1,
    32'h10F6F783,
    32'h8D3D0522,
    32'h10055533,
    32'hF37D177D,
    32'h65858082,
    32'h85934601,
    32'h06930215,
    32'hC0FB1000,
    32'h17930166,
    32'hC7B30086,
    32'h48211007,
    32'h00179713,
    32'h0007D663,
    32'h100747B3,
    32'hA0198FAD,
    32'h100747B3,
    32'h15E3187D,
    32'h112BFE08,
    32'h060500F5,
    32'h00008082,
    32'hB3B2B1B0,
    32'hB7B6B5B4,
    32'h49520001,
    32'h20564353,
    32'h2055434D,
    32'h746F6F42,
    32'h206D6F72,
    32'h50207962,
    32'h76204C43,
    32'h00302E31,
    32'h00000080,
    32'h000A3145,
    32'h0A323445,
    32'h00000000,
    32'h0A313445,
    32'h00000000,
    32'h73616C46,
    32'h44492068,
    32'h0000003A,
    32'h0A313345,
    32'h00000000,
    32'h0A323249,
    32'h00000000,
    32'h0A363245,
    32'h00000000,
    32'h43534952,
    32'h4020562D,
    32'h4C435020,
    32'h00000000,
    32'h0A323245,
    32'h00000000,
    32'h0A313245,
    32'h00000000,
    32'h0A333245,
    32'h00000000,
    32'h0A343245,
    32'h00000000,
    32'h64616F6C,
    32'h20676E69,
    32'h3A676B70,
    32'h00000000,
    32'h0A313249,
    32'h00000000,
    32'h30313245,
    32'h0000000A,
    32'h0A333249,
    32'h00000000,
    32'h0A343249,
    32'h00000000,
    32'h0A353245,
    32'h00000000,
    32'h0A373245,
    32'h00000000,
    32'h0A383245,
    32'h00000000,
    32'h0A393245,
    32'h00000000,
    32'h0A363445,
    32'h00000000,
    32'h00008D30,
    32'h00008D38,
    32'h00008D40,
    32'h00008D48,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000010,
    32'h00000000,
    32'h00527A01,
    32'h01010401,
    32'h00020D1B,
    32'h0000003C,
    32'h00000018,
    32'hFFFFF3E8,
    32'h000003A0,
    32'hC00E4200,
    32'h01115E01,
    32'h7E08117F,
    32'h117D0911,
    32'h13117C12,
    32'h7A14117B,
    32'h11791511,
    32'h17117816,
    32'h76181177,
    32'h11751911,
    32'h1B11741A,
    32'h00000073,
    32'h00000010,
    32'h00000058,
    32'hFFFFF748,
    32'h00000048,
    32'h100E4C00,
    32'h00000010,
    32'h0000006C,
    32'hFFFFF77C,
    32'h0000002C,
    32'h100E4800,
    32'h00000010,
    32'h00000080,
    32'hFFFFF794,
    32'h00000030,
    32'h00000000,
    32'h00000010,
    32'h00000094,
    32'hFFFFF7B0,
    32'h00000044,
    32'h00000000,
    32'h00000010,
    32'h000000A8,
    32'hFFFFF7E0,
    32'h00000018,
    32'h00000000,
    32'h00000010,
    32'h000000BC,
    32'hFFFFF7E4,
    32'h00000038,
    32'h100E5000,
    32'h00000010,
    32'h000000D0,
    32'hFFFFF808,
    32'h00000030,
    32'h00000000,
    32'h00000010,
    32'h000000E4,
    32'hFFFFF824,
    32'h0000001C,
    32'h100E4C00,
    32'h0000002C,
    32'h000000F8,
    32'hFFFFF82C,
    32'h0000018C,
    32'h400E4800,
    32'h7A141170,
    32'h117F0111,
    32'h09117E08,
    32'h7C12117D,
    32'h117B1311,
    32'h16117915,
    32'h77171178,
    32'h0000001C,
    32'h00000128,
    32'hFFFFF988,
    32'h0000006C,
    32'h100E4400,
    32'h7E081144,
    32'h7D09114C,
    32'h007F0111,
    32'h00000010,
    32'h00000148,
    32'hFFFFF9D4,
    32'h00000018,
    32'h00000000,
    32'h00000010,
    32'h0000015C,
    32'hFFFFF9D8,
    32'h0000005C,
    32'h00000000,
    32'h00000010,
    32'h00000170,
    32'hFFFFFA20,
    32'h0000002C,
    32'h00000000,
    32'h00000010,
    32'h00000184,
    32'hFFFFFA38,
    32'h00000024,
    32'h00000000,
    32'h00000010,
    32'h00000198,
    32'hFFFFFA48,
    32'h00000020,
    32'h00000000,
    32'h00000010,
    32'h000001AC,
    32'hFFFFFA54,
    32'h00000018,
    32'h00000000,
    32'h00000010,
    32'h000001C0,
    32'hFFFFFA58,
    32'h00000010,
    32'h00000000,
    32'h00000010,
    32'h000001D4,
    32'hFFFFFA54,
    32'h0000007C,
    32'h00000000,
    32'h0000001C,
    32'h000001E8,
    32'hFFFFFABC,
    32'h0000003E,
    32'h100E4200,
    32'h7E081146,
    32'h117D0911,
    32'h00007F01,
    32'h00000010,
    32'h00000208,
    32'hFFFFFADA,
    32'h0000001C,
    32'h00000000,
    32'h00000034,
    32'h0000021C,
    32'hFFFFFAE2,
    32'h0000018A,
    32'hC00E4200,
    32'h08114401,
    32'h7D09117E,
    32'h7C12115A,
    32'h117B1311,
    32'h01117A14,
    32'h7915117F,
    32'h11781611,
    32'h18117717,
    32'h75191176,
    32'h00000010,
    32'h00000254,
    32'hFFFFFC34,
    32'h0000002A,
    32'h00000000,
    32'h00000010,
    32'h00000268,
    32'hFFFFFC4A,
    32'h0000003C,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000};

  logic [10:0] A_Q;

  always_ff @(posedge CLK, negedge RSTN)
  begin
    if (~RSTN)
      A_Q <= '0;
    else
      if (~CSN)
        A_Q <= A;
  end

  assign Q = mem[A_Q];

endmodule